`timescale 1ns/1ps
`define DEBUG

module t_conf () ;

    reg clk ;
